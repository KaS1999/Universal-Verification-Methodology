package pack;
`include"uvm_macros.svh"
import uvm_pkg::*;
`include"seq_item.sv"
`include"sequence.sv"
`include"driver.sv"
`include"monitor.sv"
`include"agent.sv"
`include"env.sv"
`include"test.sv"
endpackage
