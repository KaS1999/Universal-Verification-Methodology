
///////////////////////////////////////PACKAGE///////////////////////////////////////////////////////
package my_package;

	`include "uvm_macros.svh"
	 import uvm_pkg::*;
     `include "seq_item.svh"
	`include "my_sequence.svh"
	`include "my_driver.svh"
	`include "my_monitor.svh"
	`include "my_agent.svh"	
	`include "my_env.svh"
	`sinclude "my_test.svh"

endpackage

